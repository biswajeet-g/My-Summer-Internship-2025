** sch_path: /home/biswajeetg/work/xschem/nmos_extract3_native.sch
**.subckt nmos_extract3_native
Vds net1 GND 1
Vsb net2 GND 0
XM3 net1 net1 net2 GND sky130_fd_pr__nfet_03v3_nvt L=0.5 W=1 nf=1 ad=0.29 as=0.29 pd=2.58 ps=2.58 nrd=0.29 nrs=0.29 sa=0 sb=0 sd=0
+ mult=1 m=1
**** begin user architecture code



.CONTROL

save all
op
write nmos_extract3_native.raw
set appendwrite
DC Vds 0 1.8 0.05 Vsb 0 0.5 0.1
write nmos_extract3_native.raw
**
plot sqrt(2*abs(Vds#branch))
plot Vds#branch

.ENDC



** opencircuitdesign pdks install
.lib /home/biswajeetg/share/pdk/sky130A/libs.tech/combined/sky130.lib.spice tt

**** end user architecture code
**.ends
.GLOBAL GND
.end
