** sch_path: /home/biswajeetg/work/xschem/nmosvds3_native.sch
**.subckt nmosvds3_native
Vgs vg GND 1
Vds vd GND 0
XM3 vd vg GND GND sky130_fd_pr__nfet_03v3_nvt L=0.5 W=1 nf=1 ad=0.29 as=0.29 pd=2.58 ps=2.58 nrd=0.29 nrs=0.29 sa=0 sb=0 sd=0
+ mult=1 m=1
**** begin user architecture code



.CONTROL

save all
OP
write nmosvds3_native.raw
set appendwrite
DC Vds 0 1.8 0.1 Vgs 0.4 1.0 0.1
write nmosvds3_native.raw
**
plot vds#branch
plot abs(vds#branch)
.ENDC



** opencircuitdesign pdks install
.lib /home/biswajeetg/share/pdk/sky130A/libs.tech/combined/sky130.lib.spice tt

**** end user architecture code
**.ends
.GLOBAL GND
.end
