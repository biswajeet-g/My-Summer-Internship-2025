** sch_path: /home/biswajeetg/work/xschem/rectifierhw.sch
**.subckt rectifierhw
V1 vin GND 0 AC 1
C1 vin vout 613f m=1
R1 vout GND 1k m=1
**** begin user architecture code



.CONTROL

save all
op
write rectifierhw.raw
set appendwrite
ac dec 10 1 10e6
write rectifierhw.raw



**** end user architecture code
**.ends
.GLOBAL GND
.end
