** sch_path: /home/biswajeetg/work/xschem/nmos_extract1.sch
**.subckt nmos_extract1
XM1 net1 net1 net2 GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1 nf=1 ad=0.29 as=0.29 pd=2.58 ps=2.58 nrd=0.29 nrs=0.29 sa=0 sb=0
+ sd=0 mult=1 m=1
Vds net1 GND 1
Vsb net2 GND 0
**** begin user architecture code



.CONTROL

save all
op
DC Vds 0 1.8 0.05 Vsb 0 0.5 0.1
plot sqrt(2*abs(Vds#branch))
plot Vds#branch

.ENDC



** opencircuitdesign pdks install
.lib /home/biswajeetg/share/pdk/sky130A/libs.tech/combined/sky130.lib.spice tt

**** end user architecture code
**.ends
.GLOBAL GND
.end
