** sch_path: /home/biswajeetg/work/xschem/currentmirrorpmos.sch
**.subckt currentmirrorpmos
Iin GND net1 50u
Vds net2 GND 1 AC 1
XM10 net2 net1 GND GND sky130_fd_pr__pfet_01v8_lvt L=1 W=4 nf=1 ad=1.16 as=1.16 pd=8.58 ps=8.58 nrd=0.0725 nrs=0.0725 sa=0 sb=0
+ sd=0 mult=1 m=1
XM1 GND net1 net1 GND sky130_fd_pr__pfet_01v8_lvt L=1 W=4 nf=1 ad=1.16 as=1.16 pd=8.58 ps=8.58 nrd=0.0725 nrs=0.0725 sa=0 sb=0
+ sd=0 mult=1 m=1
**** begin user architecture code



.CONTROL

op
write currentmirrorpmos.raw
set appendwrite
DC Vds 0 1.8 0.05
write currentmirrorpmos.raw
**
plot abs(Vds#branch)
AC dec 100 100 1000
plot '1/vm(Vds#branch)'

.ENDC




** opencircuitdesign pdks install
.lib /home/biswajeetg/share/pdk/sky130A/libs.tech/combined/sky130.lib.spice tt

**** end user architecture code
**.ends
.GLOBAL GND
.end
