** sch_path: /home/biswajeetg/work/xschem/pmos_extract1.sch
**.subckt pmos_extract1
Vds net1 GND 1
Vsb net2 GND 0
XM10 net2 net1 net1 GND sky130_fd_pr__pfet_01v8_lvt L=1 W=4 nf=1 ad=1.16 as=1.16 pd=8.58 ps=8.58 nrd=0.0725 nrs=0.0725 sa=0 sb=0
+ sd=0 mult=1 m=1
**** begin user architecture code



.CONTROL

save all
op
write pmos_extract1.raw
set appendwrite
DC Vds 0 1.8 0.05 Vsb 0 0.5 0.1
write pmos_extract1.raw
**
plot sqrt(2*abs(Vds#branch))
plot Vds#branch

.ENDC



** opencircuitdesign pdks install
.lib /home/biswajeetg/share/pdk/sky130A/libs.tech/combined/sky130.lib.spice tt

**** end user architecture code
**.ends
.GLOBAL GND
.end
